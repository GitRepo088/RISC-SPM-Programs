/*Program_Counter
*/

module Program_Counter #(
    parameter ws = 8
) (
    // count := PC_count
    output reg [ws-1: 0] count,
    // data_in := Bus_2
    input [ws-1: 0] data_in,
    input Load_PC,
    input Inc_PC,
    input clk, rst
);
    always @ (posedge clk or negedge rst)
        if(rst == 0) 
            count <= 0; 
        else if(Load_PC) 
            count <= data_in; 
        else if(Inc_PC) 
            count <= count +1;
endmodule
